
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity MUX256x8 is
	Port (
	A : 			in	std_logic_vector(255 downto 0);
	B:				out std_logic_vector(7 downto 0)
	);

end MUX256x8;

architecture Behavioral of MUX256x8 is

begin

	B <=	x"00"when A(0) = '1' else
			x"01"when A(1) = '1' else
			x"02"when A(2) = '1' else
			x"03"when A(3) = '1' else
			x"04"when A(4) = '1' else
			x"05"when A(5) = '1' else
			x"06"when A(6) = '1' else
			x"07"when A(7) = '1' else
			x"08"when A(8) = '1' else
			x"09"when A(9) = '1' else
			x"0A"when A(10) = '1' else
			x"0B"when A(11) = '1' else
			x"0C"when A(12) = '1' else
			x"0D"when A(13) = '1' else
			x"0E"when A(14) = '1' else
			x"0F"when A(15) = '1' else
			x"10"when A(16) = '1' else
			x"11"when A(17) = '1' else
			x"12"when A(18) = '1' else
			x"13"when A(19) = '1' else
			x"14"when A(20) = '1' else
			x"15"when A(21) = '1' else
			x"16"when A(22) = '1' else
			x"17"when A(23) = '1' else
			x"18"when A(24) = '1' else
			x"19"when A(25) = '1' else
			x"1A"when A(26) = '1' else
			x"1B"when A(27) = '1' else
			x"1C"when A(28) = '1' else
			x"1D"when A(29) = '1' else
			x"1E"when A(30) = '1' else
			x"1F"when A(31) = '1' else
			x"20"when A(32) = '1' else
			x"21"when A(33) = '1' else
			x"22"when A(34) = '1' else
			x"23"when A(35) = '1' else
			x"24"when A(36) = '1' else
			x"25"when A(37) = '1' else
			x"26"when A(38) = '1' else
			x"27"when A(39) = '1' else
			x"28"when A(40) = '1' else
			x"29"when A(41) = '1' else
			x"2A"when A(42) = '1' else
			x"2B"when A(43) = '1' else
			x"2C"when A(44) = '1' else
			x"2D"when A(45) = '1' else
			x"2E"when A(46) = '1' else
			x"2F"when A(47) = '1' else
			x"30"when A(48) = '1' else
			x"31"when A(49) = '1' else
			x"32"when A(50) = '1' else
			x"33"when A(51) = '1' else
			x"34"when A(52) = '1' else
			x"35"when A(53) = '1' else
			x"36"when A(54) = '1' else
			x"37"when A(55) = '1' else
			x"38"when A(56) = '1' else
			x"39"when A(57) = '1' else
			x"3A"when A(58) = '1' else
			x"3B"when A(59) = '1' else
			x"3C"when A(60) = '1' else
			x"3D"when A(61) = '1' else
			x"3E"when A(62) = '1' else
			x"3F"when A(63) = '1' else
			x"40"when A(64) = '1' else
			x"41"when A(65) = '1' else
			x"42"when A(66) = '1' else
			x"43"when A(67) = '1' else
			x"44"when A(68) = '1' else
			x"45"when A(69) = '1' else
			x"46"when A(70) = '1' else
			x"47"when A(71) = '1' else
			x"48"when A(72) = '1' else
			x"49"when A(73) = '1' else
			x"4A"when A(74) = '1' else
			x"4B"when A(75) = '1' else
			x"4C"when A(76) = '1' else
			x"4D"when A(77) = '1' else
			x"4E"when A(78) = '1' else
			x"4F"when A(79) = '1' else
			x"50"when A(80) = '1' else
			x"51"when A(81) = '1' else
			x"52"when A(82) = '1' else
			x"53"when A(83) = '1' else
			x"54"when A(84) = '1' else
			x"55"when A(85) = '1' else
			x"56"when A(86) = '1' else
			x"57"when A(87) = '1' else
			x"58"when A(88) = '1' else
			x"59"when A(89) = '1' else
			x"5A"when A(90) = '1' else
			x"5B"when A(91) = '1' else
			x"5C"when A(92) = '1' else
			x"5D"when A(93) = '1' else
			x"5E"when A(94) = '1' else
			x"5F"when A(95) = '1' else
			x"60"when A(96) = '1' else
			x"61"when A(97) = '1' else
			x"62"when A(98) = '1' else
			x"63"when A(99) = '1' else
			x"64"when A(100) = '1' else
			x"65"when A(101) = '1' else
			x"66"when A(102) = '1' else
			x"67"when A(103) = '1' else
			x"68"when A(104) = '1' else
			x"69"when A(105) = '1' else
			x"6A"when A(106) = '1' else
			x"6B"when A(107) = '1' else
			x"6C"when A(108) = '1' else
			x"6D"when A(109) = '1' else
			x"6E"when A(110) = '1' else
			x"6F"when A(111) = '1' else
			x"70"when A(112) = '1' else
			x"71"when A(113) = '1' else
			x"72"when A(114) = '1' else
			x"73"when A(115) = '1' else
			x"74"when A(116) = '1' else
			x"75"when A(117) = '1' else
			x"76"when A(118) = '1' else
			x"77"when A(119) = '1' else
			x"78"when A(120) = '1' else
			x"79"when A(121) = '1' else
			x"7A"when A(122) = '1' else
			x"7B"when A(123) = '1' else
			x"7C"when A(124) = '1' else
			x"7D"when A(125) = '1' else
			x"7E"when A(126) = '1' else
			x"7F"when A(127) = '1' else
			x"80"when A(128) = '1' else
			x"81"when A(129) = '1' else
			x"82"when A(130) = '1' else
			x"83"when A(131) = '1' else
			x"84"when A(132) = '1' else
			x"85"when A(133) = '1' else
			x"86"when A(134) = '1' else
			x"87"when A(135) = '1' else
			x"88"when A(136) = '1' else
			x"89"when A(137) = '1' else
			x"8A"when A(138) = '1' else
			x"8B"when A(139) = '1' else
			x"8C"when A(140) = '1' else
			x"8D"when A(141) = '1' else
			x"8E"when A(142) = '1' else
			x"8F"when A(143) = '1' else
			x"90"when A(144) = '1' else
			x"91"when A(145) = '1' else
			x"92"when A(146) = '1' else
			x"93"when A(147) = '1' else
			x"94"when A(148) = '1' else
			x"95"when A(149) = '1' else
			x"96"when A(150) = '1' else
			x"97"when A(151) = '1' else
			x"98"when A(152) = '1' else
			x"99"when A(153) = '1' else
			x"9A"when A(154) = '1' else
			x"9B"when A(155) = '1' else
			x"9C"when A(156) = '1' else
			x"9D"when A(157) = '1' else
			x"9E"when A(158) = '1' else
			x"9F"when A(159) = '1' else
			x"A0"when A(160) = '1' else
			x"A1"when A(161) = '1' else
			x"A2"when A(162) = '1' else
			x"A3"when A(163) = '1' else
			x"A4"when A(164) = '1' else
			x"A5"when A(165) = '1' else
			x"A6"when A(166) = '1' else
			x"A7"when A(167) = '1' else
			x"A8"when A(168) = '1' else
			x"A9"when A(169) = '1' else
			x"AA"when A(170) = '1' else
			x"AB"when A(171) = '1' else
			x"AC"when A(172) = '1' else
			x"AD"when A(173) = '1' else
			x"AE"when A(174) = '1' else
			x"AF"when A(175) = '1' else
			x"B0"when A(176) = '1' else
			x"B1"when A(177) = '1' else
			x"B2"when A(178) = '1' else
			x"B3"when A(179) = '1' else
			x"B4"when A(180) = '1' else
			x"B5"when A(181) = '1' else
			x"B6"when A(182) = '1' else
			x"B7"when A(183) = '1' else
			x"B8"when A(184) = '1' else
			x"B9"when A(185) = '1' else
			x"BA"when A(186) = '1' else
			x"BB"when A(187) = '1' else
			x"BC"when A(188) = '1' else
			x"BD"when A(189) = '1' else
			x"BE"when A(190) = '1' else
			x"BF"when A(191) = '1' else
			x"C0"when A(192) = '1' else
			x"C1"when A(193) = '1' else
			x"C2"when A(194) = '1' else
			x"C3"when A(195) = '1' else
			x"C4"when A(196) = '1' else
			x"C5"when A(197) = '1' else
			x"C6"when A(198) = '1' else
			x"C7"when A(199) = '1' else
			x"C8"when A(200) = '1' else
			x"C9"when A(201) = '1' else
			x"CA"when A(202) = '1' else
			x"CB"when A(203) = '1' else
			x"CC"when A(204) = '1' else
			x"CD"when A(205) = '1' else
			x"CE"when A(206) = '1' else
			x"CF"when A(207) = '1' else
			x"D0"when A(208) = '1' else
			x"D1"when A(209) = '1' else
			x"D2"when A(210) = '1' else
			x"D3"when A(211) = '1' else
			x"D4"when A(212) = '1' else
			x"D5"when A(213) = '1' else
			x"D6"when A(214) = '1' else
			x"D7"when A(215) = '1' else
			x"D8"when A(216) = '1' else
			x"D9"when A(217) = '1' else
			x"DA"when A(218) = '1' else
			x"DB"when A(219) = '1' else
			x"DC"when A(220) = '1' else
			x"DD"when A(221) = '1' else
			x"DE"when A(222) = '1' else
			x"DF"when A(223) = '1' else
			x"E0"when A(224) = '1' else
			x"E1"when A(225) = '1' else
			x"E2"when A(226) = '1' else
			x"E3"when A(227) = '1' else
			x"E4"when A(228) = '1' else
			x"E5"when A(229) = '1' else
			x"E6"when A(230) = '1' else
			x"E7"when A(231) = '1' else
			x"E8"when A(232) = '1' else
			x"E9"when A(233) = '1' else
			x"EA"when A(234) = '1' else
			x"EB"when A(235) = '1' else
			x"EC"when A(236) = '1' else
			x"ED"when A(237) = '1' else
			x"EE"when A(238) = '1' else
			x"EF"when A(239) = '1' else
			x"F0"when A(240) = '1' else
			x"F1"when A(241) = '1' else
			x"F2"when A(242) = '1' else
			x"F3"when A(243) = '1' else
			x"F4"when A(244) = '1' else
			x"F5"when A(245) = '1' else
			x"F6"when A(246) = '1' else
			x"F7"when A(247) = '1' else
			x"F8"when A(248) = '1' else
			x"F9"when A(249) = '1' else
			x"FA"when A(250) = '1' else
			x"FB"when A(251) = '1' else
			x"FC"when A(252) = '1' else
			x"FD"when A(253) = '1' else
			x"FE"when A(254) = '1' else
			x"FF"when A(255) = '1' else
			(others => '0');


end Behavioral;
