
-- Package for the use of AXI Stream Peripheral for Watchman
package AXIS_Peripheral_pkg is
  
  -- Register Bank Constants
	constant C_CONTROL_REG : 			integer := 0;
	constant C_NBR_OF_PACKETS_REG :		integer := 1;
	constant C_CONTENT_PACKET_1_REG :	integer := 2;
	
end AXIS_Peripheral_pkg;

package body AXIS_Peripheral_pkg is

end AXIS_Peripheral_pkg;
